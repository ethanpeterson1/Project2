library IEEE; 
use IEEE.std_logic_1164.all;
-- use work.busArray.array32;

package busArray is

type array32 is array(31 downto 0) of std_logic_vector(31 downto 0);

end package busArray;
