library IEEE;
use IEEE.std_logic_1164.all;


entity Reg_MEMWB_hw is
generic(N : integer := 137);
  port(	i_CLKn        	: in std_logic;     -- Clock input
       	i_RSTn        	: in std_logic;     -- Reset input
       	i_WEn         	: in std_logic;     -- Write enable input
	i_Flush		: in std_logic;	    -- hw

	i_ALUOut	: in std_logic_vector(31 downto 0);
	i_DMEM		: in std_logic_vector(31 downto 0);
	i_UpdatedPC	: in std_logic_vector(31 downto 0);
	i_Inst		: in std_logic_vector(31 downto 0);
	i_WriteRegAdd	: in std_logic_vector(4 downto 0);
	i_MemToReg	: in std_logic;
	i_RegWrite	: in std_logic;
	i_LuiControl	: in std_logic;
	i_JalControl	: in std_logic;

	o_ALUOut	: out std_logic_vector(31 downto 0);
	o_DMEM		: out std_logic_vector(31 downto 0);
	o_UpdatedPC	: out std_logic_vector(31 downto 0);
	o_Inst		: out std_logic_vector(31 downto 0);
	o_WriteRegAdd	: out std_logic_vector(4 downto 0);
    	o_MemToReg    	: out std_logic;
    	o_RegWrite    	: out std_logic;
	o_LuiControl	: out std_logic;
	o_JalControl	: out std_logic);

end Reg_MEMWB_hw;

architecture structural of Reg_MEMWB_hw is
component register_137 is
port(i_CLKn        : in std_logic;     -- Clock input
       i_RSTn        : in std_logic;     -- Reset input
       i_WEn         : in std_logic;     -- Write enable input
       i_Dn          : in std_logic_vector(136 downto 0);     -- Data value input
       o_Qn          : out std_logic_vector(136 downto 0));   -- Data value output
end component;

signal S_Reg_Inputs: std_logic_vector(136 downto 0);
signal S_Reg_Outputs: std_logic_vector(136 downto 0);
signal S_Flush: std_logic;					-- hw

begin
S_Reg_Inputs <= i_JalControl &
		i_LuiControl &
		i_RegWrite & 
		i_MemToReg & 
		i_WriteRegAdd &
		i_Inst &
		i_UpdatedPC &
		i_DMEM &
		i_ALUOut;

S_Flush <= i_RSTn or i_Flush;					-- hw
		
REG: register_137 port map(
	i_CLKn => i_CLKn, 
       	i_RSTn => S_Flush,					-- hw
       	i_WEn  => i_WEn,
       	i_Dn   => S_Reg_Inputs,
       	o_Qn   => S_Reg_Outputs);

o_ALUOut <= S_Reg_Outputs(31 downto 0);
o_DMEM <= S_Reg_Outputs(63 downto 32);
o_UpdatedPC <= S_Reg_Outputs(95 downto 64);
o_Inst <= S_Reg_Outputs(127 downto 96);
o_WriteRegAdd <= S_Reg_Outputs(132 downto 128);
o_MemToReg <= S_Reg_Outputs(133);
o_RegWrite <= S_Reg_Outputs(134);
o_LuiControl <= S_Reg_Outputs(135);
o_JalControl <= S_Reg_Outputs(136);


end structural;