-------------------------------------------------------------------------
-- Eduardo Contreras
-- CPR E 381
-- Lab 2
-------------------------------------------------------------------------


-- 5to32decoder.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of an edge-triggered
-- flip-flop with parallel access and reset.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity decoder5to32 is 
	port (
	      i_Sel  : in std_logic_vector(4 downto 0);
	      i_E    : in std_logic;
	      o_Dout : out std_logic_vector(31 downto 0));
	      
end decoder5to32;

architecture decoder5to32_a of decoder5to32 is
begin
   process (i_Sel, i_E)
   begin
	if (i_E = '1') then
	    case i_Sel is

		when "00000" => o_Dout <= "00000000000000000000000000000001";
		when "00001" => o_Dout <= "00000000000000000000000000000010";
		when "00010" => o_Dout <= "00000000000000000000000000000100";
		when "00011" => o_Dout <= "00000000000000000000000000001000";
		when "00100" => o_Dout <= "00000000000000000000000000010000";
		when "00101" => o_Dout <= "00000000000000000000000000100000";
		when "00110" => o_Dout <= "00000000000000000000000001000000";
		when "00111" => o_Dout <= "00000000000000000000000010000000";
		when "01000" => o_Dout <= "00000000000000000000000100000000";
		when "01001" => o_Dout <= "00000000000000000000001000000000";
		when "01010" => o_Dout <= "00000000000000000000010000000000";
		when "01011" => o_Dout <= "00000000000000000000100000000000";
		when "01100" => o_Dout <= "00000000000000000001000000000000";
		when "01101" => o_Dout <= "00000000000000000010000000000000";
		when "01110" => o_Dout <= "00000000000000000100000000000000";
		when "01111" => o_Dout <= "00000000000000001000000000000000";
		when "10000" => o_Dout <= "00000000000000010000000000000000";
		when "10001" => o_Dout <= "00000000000000100000000000000000";
		when "10010" => o_Dout <= "00000000000001000000000000000000";
		when "10011" => o_Dout <= "00000000000010000000000000000000";
		when "10100" => o_Dout <= "00000000000100000000000000000000";
		when "10101" => o_Dout <= "00000000001000000000000000000000";
		when "10110" => o_Dout <= "00000000010000000000000000000000";
		when "10111" => o_Dout <= "00000000100000000000000000000000";
		when "11000" => o_Dout <= "00000001000000000000000000000000";
		when "11001" => o_Dout <= "00000010000000000000000000000000";
		when "11010" => o_Dout <= "00000100000000000000000000000000";
		when "11011" => o_Dout <= "00001000000000000000000000000000";
		when "11100" => o_Dout <= "00010000000000000000000000000000";
		when "11101" => o_Dout <= "00100000000000000000000000000000";
		when "11110" => o_Dout <= "01000000000000000000000000000000";
		when "11111" => o_Dout <= "10000000000000000000000000000000";
		when others => o_Dout  <= "00000000000000000000000000000000";	

	    end case;
	else
		o_Dout <= "00000000000000000000000000000000";
	end if;
    end process;
end decoder5to32_a;