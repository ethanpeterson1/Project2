library IEEE;
use IEEE.std_logic_1164.all;


entity decoder32bit is

  port(i_E	: in std_logic_vector(4 downto 0);
       w_E	: in std_logic;
       o_D	: out std_logic_vector(31 downto 0));
       signal s_EnValue : std_logic_vector(5 downto 0);
end decoder32bit;

architecture dataflow of decoder32bit is
begin
	s_EnValue <= w_E & i_E;
	with s_EnValue select
		o_D <=  "00000000000000000000000000000001" when "100000",
		        "00000000000000000000000000000010" when "100001",
			"00000000000000000000000000000100" when "100010",
			"00000000000000000000000000001000" when "100011",
			"00000000000000000000000000010000" when "100100",
			"00000000000000000000000000100000" when "100101",
			"00000000000000000000000001000000" when "100110",
			"00000000000000000000000010000000" when "100111",
			"00000000000000000000000100000000" when "101000",
			"00000000000000000000001000000000" when "101001",
			"00000000000000000000010000000000" when "101010",
			"00000000000000000000100000000000" when "101011",
			"00000000000000000001000000000000" when "101100",
			"00000000000000000010000000000000" when "101101",
			"00000000000000000100000000000000" when "101110",
			"00000000000000001000000000000000" when "101111",
			"00000000000000010000000000000000" when "110000",		
			"00000000000000100000000000000000" when "110001",
			"00000000000001000000000000000000" when "110010",
			"00000000000010000000000000000000" when "110011",
			"00000000000100000000000000000000" when "110100",
			"00000000001000000000000000000000" when "110101",
			"00000000010000000000000000000000" when "110110",
			"00000000100000000000000000000000" when "110111",
			"00000001000000000000000000000000" when "111000",
			"00000010000000000000000000000000" when "111001",
			"00000100000000000000000000000000" when "111010",
			"00001000000000000000000000000000" when "111011",
			"00010000000000000000000000000000" when "111100",
			"00100000000000000000000000000000" when "111101",
			"01000000000000000000000000000000" when "111110",
			"10000000000000000000000000000000" when "111111",
			"00000000000000000000000000000000" when others;
  
end dataflow;